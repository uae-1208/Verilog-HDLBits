module top_module ( input a, input b, output out );
    mod_a m(a,b,out);
endmodule